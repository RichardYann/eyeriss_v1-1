module conv_top #(
    INWIDTH = 16
) (
    input clk,rst,
    input signed [INWIDTH-1:0]DATA_0_0
);
endmodule